module communicator(input Clk, Reset);
endmodule